module main

import client

fn main() {
	client.new_client()
}
